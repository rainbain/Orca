// Copyright 2023 Orca Hardware Emulator Project
// SPDX-License-Identifier: GPL-2.0-or-later

/*
 * RISCVSoc
 * rainbain
 * 7/4/2023
 * Orca Emulator
 *
 * XF's Top Level Logic
*/

module XFTop(
    //
    // Top Level
    //

    input wire clk, input wire resetn
);

endmodule