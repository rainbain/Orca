// Copyright 2023 Orca Hardware Emulator Project
// SPDX-License-Identifier: GPL-2.0-or-later

/*
 * WPAR
 * rainbain
 * 7/26/2023
 * Orca Emulator
 *
 * Write Gather Pipeline as used in the Gamecube.
*/

module GXFIFO(
    //
    // Top Level
    //
    input wire clk, input wire resetn,


    //
    // CPU Interface
    //
    input wire[31:0] CPUWriteData, input wire CPUWrite,


    //
    // AXI Master (Write Request Only)
    //
);

endmodule